
module gf256_power_lut (
    input [7:0] addr,
    output reg [7:0] data
);

always @(*) begin
    case(addr)
        8'd0: data = 8'h01;
        8'd1: data = 8'h03;
        8'd2: data = 8'h05;
        8'd3: data = 8'h0F;
        8'd4: data = 8'h11;
        8'd5: data = 8'h33;
        8'd6: data = 8'h55;
        8'd7: data = 8'hFF;
        8'd8: data = 8'h1A;
        8'd9: data = 8'h2E;
        8'd10: data = 8'h72;
        8'd11: data = 8'h96;
        8'd12: data = 8'hA1;
        8'd13: data = 8'hF8;
        8'd14: data = 8'h13;
        8'd15: data = 8'h35;
        8'd16: data = 8'h5F;
        8'd17: data = 8'hE1;
        8'd18: data = 8'h38;
        8'd19: data = 8'h48;
        8'd20: data = 8'hD8;
        8'd21: data = 8'h73;
        8'd22: data = 8'h95;
        8'd23: data = 8'hA4;
        8'd24: data = 8'hF7;
        8'd25: data = 8'h02;
        8'd26: data = 8'h06;
        8'd27: data = 8'h0A;
        8'd28: data = 8'h1E;
        8'd29: data = 8'h22;
        8'd30: data = 8'h66;
        8'd31: data = 8'hAA;
        8'd32: data = 8'hE5;
        8'd33: data = 8'h34;
        8'd34: data = 8'h5C;
        8'd35: data = 8'hE4;
        8'd36: data = 8'h37;
        8'd37: data = 8'h59;
        8'd38: data = 8'hEB;
        8'd39: data = 8'h26;
        8'd40: data = 8'h6A;
        8'd41: data = 8'hBE;
        8'd42: data = 8'hD9;
        8'd43: data = 8'h70;
        8'd44: data = 8'h90;
        8'd45: data = 8'hAB;
        8'd46: data = 8'hE6;
        8'd47: data = 8'h31;
        8'd48: data = 8'h53;
        8'd49: data = 8'hF5;
        8'd50: data = 8'h04;
        8'd51: data = 8'h0C;
        8'd52: data = 8'h14;
        8'd53: data = 8'h3C;
        8'd54: data = 8'h44;
        8'd55: data = 8'hCC;
        8'd56: data = 8'h4F;
        8'd57: data = 8'hD1;
        8'd58: data = 8'h68;
        8'd59: data = 8'hB8;
        8'd60: data = 8'hD3;
        8'd61: data = 8'h6E;
        8'd62: data = 8'hB2;
        8'd63: data = 8'hCD;
        8'd64: data = 8'h4C;
        8'd65: data = 8'hD4;
        8'd66: data = 8'h67;
        8'd67: data = 8'hA9;
        8'd68: data = 8'hE0;
        8'd69: data = 8'h3B;
        8'd70: data = 8'h4D;
        8'd71: data = 8'hD7;
        8'd72: data = 8'h62;
        8'd73: data = 8'hA6;
        8'd74: data = 8'hF1;
        8'd75: data = 8'h08;
        8'd76: data = 8'h18;
        8'd77: data = 8'h28;
        8'd78: data = 8'h78;
        8'd79: data = 8'h88;
        8'd80: data = 8'h83;
        8'd81: data = 8'h9E;
        8'd82: data = 8'hB9;
        8'd83: data = 8'hD0;
        8'd84: data = 8'h6B;
        8'd85: data = 8'hBD;
        8'd86: data = 8'hDC;
        8'd87: data = 8'h7F;
        8'd88: data = 8'h81;
        8'd89: data = 8'h98;
        8'd90: data = 8'hB3;
        8'd91: data = 8'hCE;
        8'd92: data = 8'h49;
        8'd93: data = 8'hDB;
        8'd94: data = 8'h76;
        8'd95: data = 8'h9A;
        8'd96: data = 8'hB5;
        8'd97: data = 8'hC4;
        8'd98: data = 8'h57;
        8'd99: data = 8'hF9;
        8'd100: data = 8'h10;
        8'd101: data = 8'h30;
        8'd102: data = 8'h50;
        8'd103: data = 8'hF0;
        8'd104: data = 8'h0B;
        8'd105: data = 8'h1D;
        8'd106: data = 8'h27;
        8'd107: data = 8'h69;
        8'd108: data = 8'hBB;
        8'd109: data = 8'hD6;
        8'd110: data = 8'h61;
        8'd111: data = 8'hA3;
        8'd112: data = 8'hFE;
        8'd113: data = 8'h19;
        8'd114: data = 8'h2B;
        8'd115: data = 8'h7D;
        8'd116: data = 8'h87;
        8'd117: data = 8'h92;
        8'd118: data = 8'hAD;
        8'd119: data = 8'hEC;
        8'd120: data = 8'h2F;
        8'd121: data = 8'h71;
        8'd122: data = 8'h93;
        8'd123: data = 8'hAE;
        8'd124: data = 8'hE9;
        8'd125: data = 8'h20;
        8'd126: data = 8'h60;
        8'd127: data = 8'hA0;
        8'd128: data = 8'hFB;
        8'd129: data = 8'h16;
        8'd130: data = 8'h3A;
        8'd131: data = 8'h4E;
        8'd132: data = 8'hD2;
        8'd133: data = 8'h6D;
        8'd134: data = 8'hB7;
        8'd135: data = 8'hC2;
        8'd136: data = 8'h5D;
        8'd137: data = 8'hE7;
        8'd138: data = 8'h32;
        8'd139: data = 8'h56;
        8'd140: data = 8'hFA;
        8'd141: data = 8'h15;
        8'd142: data = 8'h3F;
        8'd143: data = 8'h41;
        8'd144: data = 8'hC3;
        8'd145: data = 8'h5E;
        8'd146: data = 8'hE2;
        8'd147: data = 8'h3D;
        8'd148: data = 8'h47;
        8'd149: data = 8'hC9;
        8'd150: data = 8'h40;
        8'd151: data = 8'hC0;
        8'd152: data = 8'h5B;
        8'd153: data = 8'hED;
        8'd154: data = 8'h2C;
        8'd155: data = 8'h74;
        8'd156: data = 8'h9C;
        8'd157: data = 8'hBF;
        8'd158: data = 8'hDA;
        8'd159: data = 8'h75;
        8'd160: data = 8'h9F;
        8'd161: data = 8'hBA;
        8'd162: data = 8'hD5;
        8'd163: data = 8'h64;
        8'd164: data = 8'hAC;
        8'd165: data = 8'hEF;
        8'd166: data = 8'h2A;
        8'd167: data = 8'h7E;
        8'd168: data = 8'h82;
        8'd169: data = 8'h9D;
        8'd170: data = 8'hBC;
        8'd171: data = 8'hDF;
        8'd172: data = 8'h7A;
        8'd173: data = 8'h8E;
        8'd174: data = 8'h89;
        8'd175: data = 8'h80;
        8'd176: data = 8'h9B;
        8'd177: data = 8'hB6;
        8'd178: data = 8'hC1;
        8'd179: data = 8'h58;
        8'd180: data = 8'hE8;
        8'd181: data = 8'h23;
        8'd182: data = 8'h65;
        8'd183: data = 8'hAF;
        8'd184: data = 8'hEA;
        8'd185: data = 8'h25;
        8'd186: data = 8'h6F;
        8'd187: data = 8'hB1;
        8'd188: data = 8'hC8;
        8'd189: data = 8'h43;
        8'd190: data = 8'hC5;
        8'd191: data = 8'h54;
        8'd192: data = 8'hFC;
        8'd193: data = 8'h1F;
        8'd194: data = 8'h21;
        8'd195: data = 8'h63;
        8'd196: data = 8'hA5;
        8'd197: data = 8'hF4;
        8'd198: data = 8'h07;
        8'd199: data = 8'h09;
        8'd200: data = 8'h1B;
        8'd201: data = 8'h2D;
        8'd202: data = 8'h77;
        8'd203: data = 8'h99;
        8'd204: data = 8'hB0;
        8'd205: data = 8'hCB;
        8'd206: data = 8'h46;
        8'd207: data = 8'hCA;
        8'd208: data = 8'h45;
        8'd209: data = 8'hCF;
        8'd210: data = 8'h4A;
        8'd211: data = 8'hDE;
        8'd212: data = 8'h79;
        8'd213: data = 8'h8B;
        8'd214: data = 8'h86;
        8'd215: data = 8'h91;
        8'd216: data = 8'hA8;
        8'd217: data = 8'hE3;
        8'd218: data = 8'h3E;
        8'd219: data = 8'h42;
        8'd220: data = 8'hC6;
        8'd221: data = 8'h51;
        8'd222: data = 8'hF3;
        8'd223: data = 8'h0E;
        8'd224: data = 8'h12;
        8'd225: data = 8'h36;
        8'd226: data = 8'h5A;
        8'd227: data = 8'hEE;
        8'd228: data = 8'h29;
        8'd229: data = 8'h7B;
        8'd230: data = 8'h8D;
        8'd231: data = 8'h8C;
        8'd232: data = 8'h8F;
        8'd233: data = 8'h8A;
        8'd234: data = 8'h85;
        8'd235: data = 8'h94;
        8'd236: data = 8'hA7;
        8'd237: data = 8'hF2;
        8'd238: data = 8'h0D;
        8'd239: data = 8'h17;
        8'd240: data = 8'h39;
        8'd241: data = 8'h4B;
        8'd242: data = 8'hDD;
        8'd243: data = 8'h7C;
        8'd244: data = 8'h84;
        8'd245: data = 8'h97;
        8'd246: data = 8'hA2;
        8'd247: data = 8'hFD;
        8'd248: data = 8'h1C;
        8'd249: data = 8'h24;
        8'd250: data = 8'h6C;
        8'd251: data = 8'hB4;
        8'd252: data = 8'hC7;
        8'd253: data = 8'h52;
        8'd254: data = 8'hF6;
        default: data = 8'h01; // 255th power (same as 0th)
    endcase
end

endmodule
